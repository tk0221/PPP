

{-- __attribute__ syntax representation -}
nonterminal Attribute;


